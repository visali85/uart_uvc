
//This is dummy DUT. 

module dummy_dut( input clock, input reset);


endmodule

